class env;

endclass