class generator;

endclass