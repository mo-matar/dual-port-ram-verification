// Top-level testbench file that includes all components
`define WIDTH 8
`define DEPTH 256
`include "interface.sv"
`include "project_pkg.sv"
`include "../tests/basic_test.sv"
`include "tb.sv"
