// Top-level testbench file that includes all components
`include "memory_defines.sv"
`include "test_names_defines.sv"
`include "interface.sv"
`include "project_pkg.sv"
`include "basic_test.sv"
`include "write_read_tests.sv"
`include "test_factory.sv"
`include "tb.sv"
