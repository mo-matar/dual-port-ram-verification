class transaction;
endclass