class driver;




endclass