`define WIDTH 8
`define DEPTH 64
`define START_ADDR 0
`define END_ADDR (START_ADDR + `DEPTH - 1)