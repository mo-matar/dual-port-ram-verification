`define WIDTH 32
`define DEPTH 64
`define ADDR_WIDTH 16
`define START_ADDR 0
`define END_ADDR (START_ADDR + `DEPTH - 1)