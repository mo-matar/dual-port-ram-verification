// Top-level testbench file that includes all components
`include "memory_defines.sv"
`include "interface.sv"
`include "project_pkg.sv"
`include "../tests/basic_test.sv"
`include "tb.sv"
