// coverage is not needed at the moment