class scoreboard;

endclass