typedef enum {
    basic_write_read_porta,
    basic_write_read_portb,
    basic_porta_write_portb_read,
    fill_memory,
    fill_memory_porta_write_portb_read,
    fill_memory_portb_write_porta_read,
    fill_memory_porta_write_porta_read,
    fill_memory_portb_write_portb_read,
    simultaneous_read_different_address,
    simultaneous_write_different_address,
    simultaneous_write_read_same_address,
    out_of_range_memory_access,
    reset_test,
    B2B_writes_porta,
    B2B_writes_portb,
    B2B_reads_porta,
    B2B_reads_portb,
    B2B_transactions_both_ports
} test_names_e;
